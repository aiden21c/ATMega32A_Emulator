module atmega32a (
	input a,
	output b
);

assign b = a;

endmodule

