module timer_control_unit(

);

endmodule
