// Implimentation of the 8-bit Timer0 of the ATMega32A
module timer0_8bit(


);




endmodule
