module selector_32way(
	// Input selector bit
	input [4:0] S,
	
	// Output bits
	output out0,output out1,output out2,
	output out3,output out4,output out5,output out6,output out7,
	output out8,output out9,output out10,output out11,output out12,output out13,output out14,output out15,output out16,output out17,
	output out18,output out19,output out20,output out21,output out22,output out23,output out24,
	output out25,output out26,output out27,output out28,output out29,output out30,output out31
);

reg O0; reg O1; reg O2; reg O3; reg O4; reg O5; 
reg O6; reg O7; reg O8; reg O9; reg O10; reg O11; 
reg O12; reg O13; reg O14; reg O15; reg O16; reg O17; 
reg O18; reg O19; reg O20; reg O21; reg O22; reg O23; 
reg O24; reg O25; reg O26; reg O27; reg O28; reg O29; 
reg O30; reg O31; 

always @(S)
	begin
		case(S)
			5'b00000:
				begin
					O0 = 1'b1;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b00001:
				begin
					O0 = 1'b0;
					O1 = 1'b1;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b00010:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b1;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b00011:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b1;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b00100:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b1;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b00101:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b1;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b00110:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b1;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b00111:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b1;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b01000:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b1;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b01001:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b1;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b01010:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b1;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b01011:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b1;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b01100:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b1;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b01101:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b1;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b01110:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b1;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b01111:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b1;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b10000:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b1;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b10001:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b1;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b10010:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b1;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b10011:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b1;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b10100:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b1;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b10101:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b1;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b10110:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b1;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b10111:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b1;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b11000:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b1;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b11001:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b1;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b11010:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b1;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b11011:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b1;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b11100:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b1;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b11101:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b1;
					O30 = 1'b0;
					O31 = 1'b0;
				end
			5'b11110:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b1;
					O31 = 1'b0;
				end
			5'b11111:
				begin
					O0 = 1'b0;
					O1 = 1'b0;
					O2 = 1'b0;
					O3 = 1'b0;
					O4 = 1'b0;
					O5 = 1'b0;
					O6 = 1'b0;
					O7 = 1'b0;
					O8 = 1'b0;
					O9 = 1'b0;
					O10 = 1'b0;
					O11 = 1'b0;
					O12 = 1'b0;
					O13 = 1'b0;
					O14 = 1'b0;
					O15 = 1'b0;
					O16 = 1'b0;
					O17 = 1'b0;
					O18 = 1'b0;
					O19 = 1'b0;
					O20 = 1'b0;
					O21 = 1'b0;
					O22 = 1'b0;
					O23 = 1'b0;
					O24 = 1'b0;
					O25 = 1'b0;
					O26 = 1'b0;
					O27 = 1'b0;
					O28 = 1'b0;
					O29 = 1'b0;
					O30 = 1'b0;
					O31 = 1'b1;
				end
		endcase
	end



assign out0 = O0; assign out1 = O1; assign out2 = O2; assign out3 = O3; assign out4 = O4; 
assign out5 = O5; assign out6 = O6; assign out7 = O7; assign out8 = O8; assign out9 = O9; 
assign out10 = O10; assign out11 = O11; assign out12 = O12; assign out13 = O13; 
assign out14 = O14; assign out15 = O15; assign out16 = O16; assign out17 = O17; 
assign out18 = O18; assign out19 = O19; assign out20 = O20; assign out21 = O21; 
assign out22 = O22; assign out23 = O23; assign out24 = O24; assign out25 = O25; 
assign out26 = O26; assign out27 = O27; assign out28 = O28; assign out29 = O29; 
assign out30 = O30; assign out31 = O31;

endmodule
